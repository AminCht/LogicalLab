
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity multiplier is
end multiplier;

architecture Behavioral of multiplier is

begin


end Behavioral;

