
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity halfadder is
Port (
 A: in std_logic;
 B:in std_logic;
 Cin: in std_logic;
 Cout: out std_logic;
end halfadder;

architecture Behavioral of halfadder is

begin


end Behavioral;

