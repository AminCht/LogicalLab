
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity calc is
Port(
	A:in std_logic_vector(7 downto 0);
	B:in std_logic_vector(7 downto 0);
	cin:out std_logic_vector(7 downto 0));
end calc;

architecture Behavioral of calc is

begin


end Behavioral;

